`ifndef __CONFIG__
`define __CONFIG__

/*****************************************************************************/
// init file
`define MEMFILE "verification/test/test.mem"
//`define MEMFILE "verification/bench/dhrystone.mem"
//`define MEMFILE "verification/embench/wikisort.mem"
/*****************************************************************************/
// MEMORY (Byte)
`define MEM_SIZE 512*4    // 2KB (small)
//`define MEM_SIZE 1024*4   // 4KB (test)
//`define MEM_SIZE 1024*32  // 32KB (bench)
//`define MEM_SIZE 1024*64  // 64KB (embench)
/*****************************************************************************/
// start PC
`define START_PC 32'h00000000
/*****************************************************************************/
// uart queue size
`define QUEUE_SIZE 512
/*****************************************************************************/
// b = baud rate (in Mbps)
// f = frequency (in MHz) of the clk for the risc-v core (generated by clk_wiz_0)
// SERIAL_WCNT = f/b
`define SERIAL_WCNT  40   // default 100
/*****************************************************************************/

`endif
